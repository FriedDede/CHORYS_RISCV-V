/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
// 21/03/2025 10:31:48
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o,
   output logic         rvalid_o
);
    localparam int RomSize = 408;

    const logic [RomSize-1:0][63:0] mem = {
        64'h0000040c_00000400,
        64'h000003f4_000003e8,
        64'h000003dc_000003d0,
        64'h000003c4_000003b8,
        64'h000003ac_000003a0,
        64'h00000394_00000388,
        64'h0000037c_00000370,
        64'h00000364_00000358,
        64'h0000034c_00000340,
        64'h00000334_00000328,
        64'h0000031c_00000310,
        64'h00000304_000002f4,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hee9ff06f_000400e7,
        64'h97010437_ef5ff06f,
        64'h000400e7_96010437,
        64'hf01ff06f_000400e7,
        64'h95010437_f0dff06f,
        64'h000400e7_94010437,
        64'hf19ff06f_000400e7,
        64'h93010437_f25ff06f,
        64'h000400e7_92010437,
        64'hf31ff06f_000400e7,
        64'h91010437_f3dff06f,
        64'h000400e7_90010437,
        64'hf49ff06f_000400e7,
        64'h8f010437_f55ff06f,
        64'h000400e7_8e010437,
        64'hf61ff06f_000400e7,
        64'h8d010437_f6dff06f,
        64'h000400e7_8c010437,
        64'hf79ff06f_000400e7,
        64'h8b010437_f85ff06f,
        64'h000400e7_8a010437,
        64'hf91ff06f_000400e7,
        64'h89010437_f9dff06f,
        64'h000400e7_88010437,
        64'hfa9ff06f_000400e7,
        64'h87010437_fb5ff06f,
        64'h000400e7_86010437,
        64'hfc1ff06f_000400e7,
        64'h85010437_fcdff06f,
        64'h000400e7_84010437,
        64'hfd9ff06f_000400e7,
        64'h83010437_fe5ff06f,
        64'h000400e7_82010437,
        64'hff1ff06f_000400e7,
        64'h81010437_00008067,
        64'h00000513_000400e7,
        64'h80010437_00078067,
        64'h0007a783_00e787b3,
        64'h60000713_00279793,
        64'h02f76063_01700713,
        64'hf14027f3_e55ff06f,
        64'h02010113_01c12083,
        64'h00d14503_e65ff0ef,
        64'h00c14503_f0dff0ef,
        64'h00112e23_00c10593,
        64'hfe010113_00008067,
        64'h02010113_01012903,
        64'h01412483_01812403,
        64'h01c12083_fd241ee3,
        64'he99ff0ef_00d14503,
        64'hea1ff0ef_ff840413,
        64'h00c14503_f4dff0ef,
        64'h0ff57513_00c10593,
        64'h0084d533_ff800913,
        64'h03800413_00050493,
        64'h00112e23_01212823,
        64'h00912a23_00812c23,
        64'hfe010113_00008067,
        64'h02010113_01012903,
        64'h01412483_01812403,
        64'h01c12083_fd241ee3,
        64'hef9ff0ef_00d14503,
        64'hf01ff0ef_ff840413,
        64'h00c14503_fadff0ef,
        64'h0ff57513_00c10593,
        64'h0084d533_ff800913,
        64'h01800413_00050493,
        64'h00112e23_01212823,
        64'h00912a23_00812c23,
        64'hfe010113_00008067,
        64'h00f58023_0007c783,
        64'h00e580a3_00a787b3,
        64'h00455513_00074703,
        64'h00e78733_00f57713,
        64'h50000793_fe1ff06f,
        64'h00140413_f6dff0ef,
        64'h00008067_01010113,
        64'h00812403_00c12083,
        64'h00051a63_00044503,
        64'h00050413_00112623,
        64'h00812423_ff010113,
        64'h00008067_00e78823,
        64'h02000713_00e78423,
        64'hfc700713_00e78623,
        64'h00300713_00a70223,
        64'h0ff57513_00c70023,
        64'h00855513_0ff57613,
        64'h00070793_00d70623,
        64'hf8000693_00070223,
        64'h14000737_02b55533,
        64'h00459593_00008067,
        64'h00a78023_140007b7,
        64'hfe078ce3_0207f793,
        64'h00074783_01470713,
        64'h14000737_00008067,
        64'h02057513_0147c503,
        64'h140007b7_00008067,
        64'h00054503_00008067,
        64'h00b50023_0000006f,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000006f_2bc000ef,
        64'h90000137_30029073,
        64'h000022b7_30529073,
        64'h10028293_00000297
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
            rvalid_o <= 1;
        end else begin
            rvalid_o <= 0;
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
